module top;

   bit clk, rst_n;

   clock_unit clock(clk);
   test test();

endmodule
