module bindfiles;
   bind dut dut_asserts p1 (.*);
endmodule
